module onehot_tb #(
	parameter int W = 4,
	parameter bit MSB = 1
)
(
	input wire [W-1:0] i,
	output reg [W-1:0] o
);

endmodule
